module main;
  initial
    begin
      $display("Fuck You Github!");
      $finish;
    end
endmodule
